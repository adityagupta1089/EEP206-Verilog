module full_adder (a,b,cin,s,cout);
  input a,b,cin;
  output s,cout;
  assign s=a^b^cin;
  assign cout=(a&b)|(b&cin)|(cin&a);
endmodule // full_adder
module four_bit_ripple_adder (a,b,sum,cout);
  input [3:0] a,b;
  wire [2:0] c;
  output [3:0] sum;
  output cout;
  full_adder fa1(a[0],b[0],0,sum[0],c[0]);
  full_adder fa2(a[1],b[1],c[0],sum[1],c[1]);
  full_adder fa3(a[2],b[2],c[1],sum[2],c[2]);
  full_adder fa4(a[3],b[3],c[2],sum[3],cout);
endmodule // 4_bit_ripple_adder
module four_bit_ripple_adder_tb;

reg [3:0] a,b;
wire [3:0] s;
wire c;

four_bit_ripple_adder fbra (.a(a),.b(b),.sum(s),.cout(c));

initial begin
  $monitor ("a=%b, b=%b, s=%b, c=%b",a,b,s,c);
  a=4'b0; b=4'b0;
#5 a=4'b0; b=4'b1;
#5 a=4'b0; b=4'b10;
#5 a=4'b0; b=4'b11;
#5 a=4'b0; b=4'b100;
#5 a=4'b0; b=4'b101;
#5 a=4'b0; b=4'b110;
#5 a=4'b0; b=4'b111;
#5 a=4'b0; b=4'b1000;
#5 a=4'b0; b=4'b1001;
#5 a=4'b0; b=4'b1010;
#5 a=4'b0; b=4'b1011;
#5 a=4'b0; b=4'b1100;
#5 a=4'b0; b=4'b1101;
#5 a=4'b0; b=4'b1110;
#5 a=4'b0; b=4'b1111;
#5 a=4'b1; b=4'b0;
#5 a=4'b1; b=4'b1;
#5 a=4'b1; b=4'b10;
#5 a=4'b1; b=4'b11;
#5 a=4'b1; b=4'b100;
#5 a=4'b1; b=4'b101;
#5 a=4'b1; b=4'b110;
#5 a=4'b1; b=4'b111;
#5 a=4'b1; b=4'b1000;
#5 a=4'b1; b=4'b1001;
#5 a=4'b1; b=4'b1010;
#5 a=4'b1; b=4'b1011;
#5 a=4'b1; b=4'b1100;
#5 a=4'b1; b=4'b1101;
#5 a=4'b1; b=4'b1110;
#5 a=4'b1; b=4'b1111;
#5 a=4'b10; b=4'b0;
#5 a=4'b10; b=4'b1;
#5 a=4'b10; b=4'b10;
#5 a=4'b10; b=4'b11;
#5 a=4'b10; b=4'b100;
#5 a=4'b10; b=4'b101;
#5 a=4'b10; b=4'b110;
#5 a=4'b10; b=4'b111;
#5 a=4'b10; b=4'b1000;
#5 a=4'b10; b=4'b1001;
#5 a=4'b10; b=4'b1010;
#5 a=4'b10; b=4'b1011;
#5 a=4'b10; b=4'b1100;
#5 a=4'b10; b=4'b1101;
#5 a=4'b10; b=4'b1110;
#5 a=4'b10; b=4'b1111;
#5 a=4'b11; b=4'b0;
#5 a=4'b11; b=4'b1;
#5 a=4'b11; b=4'b10;
#5 a=4'b11; b=4'b11;
#5 a=4'b11; b=4'b100;
#5 a=4'b11; b=4'b101;
#5 a=4'b11; b=4'b110;
#5 a=4'b11; b=4'b111;
#5 a=4'b11; b=4'b1000;
#5 a=4'b11; b=4'b1001;
#5 a=4'b11; b=4'b1010;
#5 a=4'b11; b=4'b1011;
#5 a=4'b11; b=4'b1100;
#5 a=4'b11; b=4'b1101;
#5 a=4'b11; b=4'b1110;
#5 a=4'b11; b=4'b1111;
#5 a=4'b100; b=4'b0;
#5 a=4'b100; b=4'b1;
#5 a=4'b100; b=4'b10;
#5 a=4'b100; b=4'b11;
#5 a=4'b100; b=4'b100;
#5 a=4'b100; b=4'b101;
#5 a=4'b100; b=4'b110;
#5 a=4'b100; b=4'b111;
#5 a=4'b100; b=4'b1000;
#5 a=4'b100; b=4'b1001;
#5 a=4'b100; b=4'b1010;
#5 a=4'b100; b=4'b1011;
#5 a=4'b100; b=4'b1100;
#5 a=4'b100; b=4'b1101;
#5 a=4'b100; b=4'b1110;
#5 a=4'b100; b=4'b1111;
#5 a=4'b101; b=4'b0;
#5 a=4'b101; b=4'b1;
#5 a=4'b101; b=4'b10;
#5 a=4'b101; b=4'b11;
#5 a=4'b101; b=4'b100;
#5 a=4'b101; b=4'b101;
#5 a=4'b101; b=4'b110;
#5 a=4'b101; b=4'b111;
#5 a=4'b101; b=4'b1000;
#5 a=4'b101; b=4'b1001;
#5 a=4'b101; b=4'b1010;
#5 a=4'b101; b=4'b1011;
#5 a=4'b101; b=4'b1100;
#5 a=4'b101; b=4'b1101;
#5 a=4'b101; b=4'b1110;
#5 a=4'b101; b=4'b1111;
#5 a=4'b110; b=4'b0;
#5 a=4'b110; b=4'b1;
#5 a=4'b110; b=4'b10;
#5 a=4'b110; b=4'b11;
#5 a=4'b110; b=4'b100;
#5 a=4'b110; b=4'b101;
#5 a=4'b110; b=4'b110;
#5 a=4'b110; b=4'b111;
#5 a=4'b110; b=4'b1000;
#5 a=4'b110; b=4'b1001;
#5 a=4'b110; b=4'b1010;
#5 a=4'b110; b=4'b1011;
#5 a=4'b110; b=4'b1100;
#5 a=4'b110; b=4'b1101;
#5 a=4'b110; b=4'b1110;
#5 a=4'b110; b=4'b1111;
#5 a=4'b111; b=4'b0;
#5 a=4'b111; b=4'b1;
#5 a=4'b111; b=4'b10;
#5 a=4'b111; b=4'b11;
#5 a=4'b111; b=4'b100;
#5 a=4'b111; b=4'b101;
#5 a=4'b111; b=4'b110;
#5 a=4'b111; b=4'b111;
#5 a=4'b111; b=4'b1000;
#5 a=4'b111; b=4'b1001;
#5 a=4'b111; b=4'b1010;
#5 a=4'b111; b=4'b1011;
#5 a=4'b111; b=4'b1100;
#5 a=4'b111; b=4'b1101;
#5 a=4'b111; b=4'b1110;
#5 a=4'b111; b=4'b1111;
#5 a=4'b1000; b=4'b0;
#5 a=4'b1000; b=4'b1;
#5 a=4'b1000; b=4'b10;
#5 a=4'b1000; b=4'b11;
#5 a=4'b1000; b=4'b100;
#5 a=4'b1000; b=4'b101;
#5 a=4'b1000; b=4'b110;
#5 a=4'b1000; b=4'b111;
#5 a=4'b1000; b=4'b1000;
#5 a=4'b1000; b=4'b1001;
#5 a=4'b1000; b=4'b1010;
#5 a=4'b1000; b=4'b1011;
#5 a=4'b1000; b=4'b1100;
#5 a=4'b1000; b=4'b1101;
#5 a=4'b1000; b=4'b1110;
#5 a=4'b1000; b=4'b1111;
#5 a=4'b1001; b=4'b0;
#5 a=4'b1001; b=4'b1;
#5 a=4'b1001; b=4'b10;
#5 a=4'b1001; b=4'b11;
#5 a=4'b1001; b=4'b100;
#5 a=4'b1001; b=4'b101;
#5 a=4'b1001; b=4'b110;
#5 a=4'b1001; b=4'b111;
#5 a=4'b1001; b=4'b1000;
#5 a=4'b1001; b=4'b1001;
#5 a=4'b1001; b=4'b1010;
#5 a=4'b1001; b=4'b1011;
#5 a=4'b1001; b=4'b1100;
#5 a=4'b1001; b=4'b1101;
#5 a=4'b1001; b=4'b1110;
#5 a=4'b1001; b=4'b1111;
#5 a=4'b1010; b=4'b0;
#5 a=4'b1010; b=4'b1;
#5 a=4'b1010; b=4'b10;
#5 a=4'b1010; b=4'b11;
#5 a=4'b1010; b=4'b100;
#5 a=4'b1010; b=4'b101;
#5 a=4'b1010; b=4'b110;
#5 a=4'b1010; b=4'b111;
#5 a=4'b1010; b=4'b1000;
#5 a=4'b1010; b=4'b1001;
#5 a=4'b1010; b=4'b1010;
#5 a=4'b1010; b=4'b1011;
#5 a=4'b1010; b=4'b1100;
#5 a=4'b1010; b=4'b1101;
#5 a=4'b1010; b=4'b1110;
#5 a=4'b1010; b=4'b1111;
#5 a=4'b1011; b=4'b0;
#5 a=4'b1011; b=4'b1;
#5 a=4'b1011; b=4'b10;
#5 a=4'b1011; b=4'b11;
#5 a=4'b1011; b=4'b100;
#5 a=4'b1011; b=4'b101;
#5 a=4'b1011; b=4'b110;
#5 a=4'b1011; b=4'b111;
#5 a=4'b1011; b=4'b1000;
#5 a=4'b1011; b=4'b1001;
#5 a=4'b1011; b=4'b1010;
#5 a=4'b1011; b=4'b1011;
#5 a=4'b1011; b=4'b1100;
#5 a=4'b1011; b=4'b1101;
#5 a=4'b1011; b=4'b1110;
#5 a=4'b1011; b=4'b1111;
#5 a=4'b1100; b=4'b0;
#5 a=4'b1100; b=4'b1;
#5 a=4'b1100; b=4'b10;
#5 a=4'b1100; b=4'b11;
#5 a=4'b1100; b=4'b100;
#5 a=4'b1100; b=4'b101;
#5 a=4'b1100; b=4'b110;
#5 a=4'b1100; b=4'b111;
#5 a=4'b1100; b=4'b1000;
#5 a=4'b1100; b=4'b1001;
#5 a=4'b1100; b=4'b1010;
#5 a=4'b1100; b=4'b1011;
#5 a=4'b1100; b=4'b1100;
#5 a=4'b1100; b=4'b1101;
#5 a=4'b1100; b=4'b1110;
#5 a=4'b1100; b=4'b1111;
#5 a=4'b1101; b=4'b0;
#5 a=4'b1101; b=4'b1;
#5 a=4'b1101; b=4'b10;
#5 a=4'b1101; b=4'b11;
#5 a=4'b1101; b=4'b100;
#5 a=4'b1101; b=4'b101;
#5 a=4'b1101; b=4'b110;
#5 a=4'b1101; b=4'b111;
#5 a=4'b1101; b=4'b1000;
#5 a=4'b1101; b=4'b1001;
#5 a=4'b1101; b=4'b1010;
#5 a=4'b1101; b=4'b1011;
#5 a=4'b1101; b=4'b1100;
#5 a=4'b1101; b=4'b1101;
#5 a=4'b1101; b=4'b1110;
#5 a=4'b1101; b=4'b1111;
#5 a=4'b1110; b=4'b0;
#5 a=4'b1110; b=4'b1;
#5 a=4'b1110; b=4'b10;
#5 a=4'b1110; b=4'b11;
#5 a=4'b1110; b=4'b100;
#5 a=4'b1110; b=4'b101;
#5 a=4'b1110; b=4'b110;
#5 a=4'b1110; b=4'b111;
#5 a=4'b1110; b=4'b1000;
#5 a=4'b1110; b=4'b1001;
#5 a=4'b1110; b=4'b1010;
#5 a=4'b1110; b=4'b1011;
#5 a=4'b1110; b=4'b1100;
#5 a=4'b1110; b=4'b1101;
#5 a=4'b1110; b=4'b1110;
#5 a=4'b1110; b=4'b1111;
#5 a=4'b1111; b=4'b0;
#5 a=4'b1111; b=4'b1;
#5 a=4'b1111; b=4'b10;
#5 a=4'b1111; b=4'b11;
#5 a=4'b1111; b=4'b100;
#5 a=4'b1111; b=4'b101;
#5 a=4'b1111; b=4'b110;
#5 a=4'b1111; b=4'b111;
#5 a=4'b1111; b=4'b1000;
#5 a=4'b1111; b=4'b1001;
#5 a=4'b1111; b=4'b1010;
#5 a=4'b1111; b=4'b1011;
#5 a=4'b1111; b=4'b1100;
#5 a=4'b1111; b=4'b1101;
#5 a=4'b1111; b=4'b1110;
#5 a=4'b1111; b=4'b1111;
  $finish;
end

endmodule // four_bit_ripple_adder_tb

/*Output:
a=0000, b=0000, s=0000, c=0
a=0000, b=0001, s=0001, c=0
a=0000, b=0010, s=0010, c=0
a=0000, b=0011, s=0011, c=0
a=0000, b=0100, s=0100, c=0
a=0000, b=0101, s=0101, c=0
a=0000, b=0110, s=0110, c=0
a=0000, b=0111, s=0111, c=0
a=0000, b=1000, s=1000, c=0
a=0000, b=1001, s=1001, c=0
a=0000, b=1010, s=1010, c=0
a=0000, b=1011, s=1011, c=0
a=0000, b=1100, s=1100, c=0
a=0000, b=1101, s=1101, c=0
a=0000, b=1110, s=1110, c=0
a=0000, b=1111, s=1111, c=0
a=0001, b=0000, s=0001, c=0
a=0001, b=0001, s=0010, c=0
a=0001, b=0010, s=0011, c=0
a=0001, b=0011, s=0100, c=0
a=0001, b=0100, s=0101, c=0
a=0001, b=0101, s=0110, c=0
a=0001, b=0110, s=0111, c=0
a=0001, b=0111, s=1000, c=0
a=0001, b=1000, s=1001, c=0
a=0001, b=1001, s=1010, c=0
a=0001, b=1010, s=1011, c=0
a=0001, b=1011, s=1100, c=0
a=0001, b=1100, s=1101, c=0
a=0001, b=1101, s=1110, c=0
a=0001, b=1110, s=1111, c=0
a=0001, b=1111, s=0000, c=1
a=0010, b=0000, s=0010, c=0
a=0010, b=0001, s=0011, c=0
a=0010, b=0010, s=0100, c=0
a=0010, b=0011, s=0101, c=0
a=0010, b=0100, s=0110, c=0
a=0010, b=0101, s=0111, c=0
a=0010, b=0110, s=1000, c=0
a=0010, b=0111, s=1001, c=0
a=0010, b=1000, s=1010, c=0
a=0010, b=1001, s=1011, c=0
a=0010, b=1010, s=1100, c=0
a=0010, b=1011, s=1101, c=0
a=0010, b=1100, s=1110, c=0
a=0010, b=1101, s=1111, c=0
a=0010, b=1110, s=0000, c=1
a=0010, b=1111, s=0001, c=1
a=0011, b=0000, s=0011, c=0
a=0011, b=0001, s=0100, c=0
a=0011, b=0010, s=0101, c=0
a=0011, b=0011, s=0110, c=0
a=0011, b=0100, s=0111, c=0
a=0011, b=0101, s=1000, c=0
a=0011, b=0110, s=1001, c=0
a=0011, b=0111, s=1010, c=0
a=0011, b=1000, s=1011, c=0
a=0011, b=1001, s=1100, c=0
a=0011, b=1010, s=1101, c=0
a=0011, b=1011, s=1110, c=0
a=0011, b=1100, s=1111, c=0
a=0011, b=1101, s=0000, c=1
a=0011, b=1110, s=0001, c=1
a=0011, b=1111, s=0010, c=1
a=0100, b=0000, s=0100, c=0
a=0100, b=0001, s=0101, c=0
a=0100, b=0010, s=0110, c=0
a=0100, b=0011, s=0111, c=0
a=0100, b=0100, s=1000, c=0
a=0100, b=0101, s=1001, c=0
a=0100, b=0110, s=1010, c=0
a=0100, b=0111, s=1011, c=0
a=0100, b=1000, s=1100, c=0
a=0100, b=1001, s=1101, c=0
a=0100, b=1010, s=1110, c=0
a=0100, b=1011, s=1111, c=0
a=0100, b=1100, s=0000, c=1
a=0100, b=1101, s=0001, c=1
a=0100, b=1110, s=0010, c=1
a=0100, b=1111, s=0011, c=1
a=0101, b=0000, s=0101, c=0
a=0101, b=0001, s=0110, c=0
a=0101, b=0010, s=0111, c=0
a=0101, b=0011, s=1000, c=0
a=0101, b=0100, s=1001, c=0
a=0101, b=0101, s=1010, c=0
a=0101, b=0110, s=1011, c=0
a=0101, b=0111, s=1100, c=0
a=0101, b=1000, s=1101, c=0
a=0101, b=1001, s=1110, c=0
a=0101, b=1010, s=1111, c=0
a=0101, b=1011, s=0000, c=1
a=0101, b=1100, s=0001, c=1
a=0101, b=1101, s=0010, c=1
a=0101, b=1110, s=0011, c=1
a=0101, b=1111, s=0100, c=1
a=0110, b=0000, s=0110, c=0
a=0110, b=0001, s=0111, c=0
a=0110, b=0010, s=1000, c=0
a=0110, b=0011, s=1001, c=0
a=0110, b=0100, s=1010, c=0
a=0110, b=0101, s=1011, c=0
a=0110, b=0110, s=1100, c=0
a=0110, b=0111, s=1101, c=0
a=0110, b=1000, s=1110, c=0
a=0110, b=1001, s=1111, c=0
a=0110, b=1010, s=0000, c=1
a=0110, b=1011, s=0001, c=1
a=0110, b=1100, s=0010, c=1
a=0110, b=1101, s=0011, c=1
a=0110, b=1110, s=0100, c=1
a=0110, b=1111, s=0101, c=1
a=0111, b=0000, s=0111, c=0
a=0111, b=0001, s=1000, c=0
a=0111, b=0010, s=1001, c=0
a=0111, b=0011, s=1010, c=0
a=0111, b=0100, s=1011, c=0
a=0111, b=0101, s=1100, c=0
a=0111, b=0110, s=1101, c=0
a=0111, b=0111, s=1110, c=0
a=0111, b=1000, s=1111, c=0
a=0111, b=1001, s=0000, c=1
a=0111, b=1010, s=0001, c=1
a=0111, b=1011, s=0010, c=1
a=0111, b=1100, s=0011, c=1
a=0111, b=1101, s=0100, c=1
a=0111, b=1110, s=0101, c=1
a=0111, b=1111, s=0110, c=1
a=1000, b=0000, s=1000, c=0
a=1000, b=0001, s=1001, c=0
a=1000, b=0010, s=1010, c=0
a=1000, b=0011, s=1011, c=0
a=1000, b=0100, s=1100, c=0
a=1000, b=0101, s=1101, c=0
a=1000, b=0110, s=1110, c=0
a=1000, b=0111, s=1111, c=0
a=1000, b=1000, s=0000, c=1
a=1000, b=1001, s=0001, c=1
a=1000, b=1010, s=0010, c=1
a=1000, b=1011, s=0011, c=1
a=1000, b=1100, s=0100, c=1
a=1000, b=1101, s=0101, c=1
a=1000, b=1110, s=0110, c=1
a=1000, b=1111, s=0111, c=1
a=1001, b=0000, s=1001, c=0
a=1001, b=0001, s=1010, c=0
a=1001, b=0010, s=1011, c=0
a=1001, b=0011, s=1100, c=0
a=1001, b=0100, s=1101, c=0
a=1001, b=0101, s=1110, c=0
a=1001, b=0110, s=1111, c=0
a=1001, b=0111, s=0000, c=1
a=1001, b=1000, s=0001, c=1
a=1001, b=1001, s=0010, c=1
a=1001, b=1010, s=0011, c=1
a=1001, b=1011, s=0100, c=1
a=1001, b=1100, s=0101, c=1
a=1001, b=1101, s=0110, c=1
a=1001, b=1110, s=0111, c=1
a=1001, b=1111, s=1000, c=1
a=1010, b=0000, s=1010, c=0
a=1010, b=0001, s=1011, c=0
a=1010, b=0010, s=1100, c=0
a=1010, b=0011, s=1101, c=0
a=1010, b=0100, s=1110, c=0
a=1010, b=0101, s=1111, c=0
a=1010, b=0110, s=0000, c=1
a=1010, b=0111, s=0001, c=1
a=1010, b=1000, s=0010, c=1
a=1010, b=1001, s=0011, c=1
a=1010, b=1010, s=0100, c=1
a=1010, b=1011, s=0101, c=1
a=1010, b=1100, s=0110, c=1
a=1010, b=1101, s=0111, c=1
a=1010, b=1110, s=1000, c=1
a=1010, b=1111, s=1001, c=1
a=1011, b=0000, s=1011, c=0
a=1011, b=0001, s=1100, c=0
a=1011, b=0010, s=1101, c=0
a=1011, b=0011, s=1110, c=0
a=1011, b=0100, s=1111, c=0
a=1011, b=0101, s=0000, c=1
a=1011, b=0110, s=0001, c=1
a=1011, b=0111, s=0010, c=1
a=1011, b=1000, s=0011, c=1
a=1011, b=1001, s=0100, c=1
a=1011, b=1010, s=0101, c=1
a=1011, b=1011, s=0110, c=1
a=1011, b=1100, s=0111, c=1
a=1011, b=1101, s=1000, c=1
a=1011, b=1110, s=1001, c=1
a=1011, b=1111, s=1010, c=1
a=1100, b=0000, s=1100, c=0
a=1100, b=0001, s=1101, c=0
a=1100, b=0010, s=1110, c=0
a=1100, b=0011, s=1111, c=0
a=1100, b=0100, s=0000, c=1
a=1100, b=0101, s=0001, c=1
a=1100, b=0110, s=0010, c=1
a=1100, b=0111, s=0011, c=1
a=1100, b=1000, s=0100, c=1
a=1100, b=1001, s=0101, c=1
a=1100, b=1010, s=0110, c=1
a=1100, b=1011, s=0111, c=1
a=1100, b=1100, s=1000, c=1
a=1100, b=1101, s=1001, c=1
a=1100, b=1110, s=1010, c=1
a=1100, b=1111, s=1011, c=1
a=1101, b=0000, s=1101, c=0
a=1101, b=0001, s=1110, c=0
a=1101, b=0010, s=1111, c=0
a=1101, b=0011, s=0000, c=1
a=1101, b=0100, s=0001, c=1
a=1101, b=0101, s=0010, c=1
a=1101, b=0110, s=0011, c=1
a=1101, b=0111, s=0100, c=1
a=1101, b=1000, s=0101, c=1
a=1101, b=1001, s=0110, c=1
a=1101, b=1010, s=0111, c=1
a=1101, b=1011, s=1000, c=1
a=1101, b=1100, s=1001, c=1
a=1101, b=1101, s=1010, c=1
a=1101, b=1110, s=1011, c=1
a=1101, b=1111, s=1100, c=1
a=1110, b=0000, s=1110, c=0
a=1110, b=0001, s=1111, c=0
a=1110, b=0010, s=0000, c=1
a=1110, b=0011, s=0001, c=1
a=1110, b=0100, s=0010, c=1
a=1110, b=0101, s=0011, c=1
a=1110, b=0110, s=0100, c=1
a=1110, b=0111, s=0101, c=1
a=1110, b=1000, s=0110, c=1
a=1110, b=1001, s=0111, c=1
a=1110, b=1010, s=1000, c=1
a=1110, b=1011, s=1001, c=1
a=1110, b=1100, s=1010, c=1
a=1110, b=1101, s=1011, c=1
a=1110, b=1110, s=1100, c=1
a=1110, b=1111, s=1101, c=1
a=1111, b=0000, s=1111, c=0
a=1111, b=0001, s=0000, c=1
a=1111, b=0010, s=0001, c=1
a=1111, b=0011, s=0010, c=1
a=1111, b=0100, s=0011, c=1
a=1111, b=0101, s=0100, c=1
a=1111, b=0110, s=0101, c=1
a=1111, b=0111, s=0110, c=1
a=1111, b=1000, s=0111, c=1
a=1111, b=1001, s=1000, c=1
a=1111, b=1010, s=1001, c=1
a=1111, b=1011, s=1010, c=1
a=1111, b=1100, s=1011, c=1
a=1111, b=1101, s=1100, c=1
a=1111, b=1110, s=1101, c=1
a=1111, b=1111, s=1110, c=1
*/
